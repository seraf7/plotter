library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_ARITH.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;


entity octagono is
	 generic( Max: natural := 1000000);
    Port ( reloj : in  STD_LOGIC;
			  inicio: in STD_LOGIC;
			  movServo : out STD_LOGIC;
			  En0, En1, dir0, dir1 : out STD_LOGIC
         );
end octagono;

architecture Behavioral of octagono is

signal PWM_Count: integer range 1 to Max;--1000000;

signal seg, selector: std_logic;
signal cont: integer;


--Biblioteca de estados
type Estados is (S0, S1, S2, S3, S4, S5, S6, S7, S8, S9);
signal epresente, esiguiente: Estados;

begin

generacion_PWM: process(reloj, selector, PWM_Count)
    constant pos1: integer := 50000;  --representa a 1.00ms = 0°
    constant pos4: integer := 100000; --representa a 2.00ms = 180°
        begin
        if rising_edge(reloj) then 
            PWM_Count <= PWM_Count + 1;
        end if;
        case (selector) is
            when '1' =>--con el selector en 1 se posiciona en servo en 0°
                if PWM_Count <= pos1 then
                    movServo <= '1';
                else
                    movServo <= '0';
                end if;
            when others =>-- con el selector en 0 se posiciona en servo en 180°
                if PWM_Count <= pos4 then
                    movServo <= '1';
                else
                    movServo <= '0';
                end if;
        end case;
    end process generacion_PWM;

-----------
	divi: process(reloj)
	variable toggle: std_logic:='0';
	variable cuenta: std_logic_vector(27 downto 0):=X"0000000";		--Declaracion de una varible interna de proceso
	begin
		if rising_edge (reloj) then
			if cuenta = X"003D090" then		--Tiempo para 0.5s,  2BA3487,   04C4B40
				toggle := NOT(toggle); 
				cuenta:=X"0000000";
			else
				cuenta:= cuenta + 1;
			end if;
		end if;
		seg <= toggle; ---modificacion de frecuencia
	end process;
	
ASM1: process(seg)
variable cuenta:  integer := 0;
begin
	if rising_edge(seg) then
		if epresente = esiguiente then 
			cuenta:=cuenta+1;
		else
			cuenta:= 0;
		end if;
		epresente <= esiguiente;
	end if;
cont<=cuenta;
end process;

ASM2: process(epresente,cont)

begin

	case epresente is
		when S0 =>
			selector <= '1';
			En0 <= '0';
			En1 <= '0';
			dir0 <= '0';
			dir1 <= '0';
			if inicio = '1' then
				esiguiente<= S1;
				selector <= '0';
			else
				esiguiente <= S0;
			end if;
			
		when S1 =>
			selector <= '0';
			En0 <= '0';
			En1 <= '0';
			dir0 <= '1';
			dir1 <= '0';	
			esiguiente <= S2;
		
		when S2 =>
			selector <= '0';
			En0 <= '1';
			En1 <= '0';
			dir0 <= '1';
			dir1 <= '1';
			if cont = 250 then --Contamos hasta 15, 340
				esiguiente<=S3;
			else
				esiguiente<=S2;
			end if;
		
		when S3 =>
			selector <= '0';
			En0 <= '1';
			En1 <= '1';
			dir0 <= '1';
			dir1 <= '1';
			if cont = 133 then --Contamos hasta 15, 340
				esiguiente<=S4;
			else
				esiguiente<=S3;
			end if;
			
		when S4 =>
			selector <= '0';
			En0 <= '0';
			En1 <= '1';
			dir0 <= '0';
			dir1 <= '1';
			if cont = 250 then --Contamos hasta 15
				esiguiente<=S5;
			else
				esiguiente<=S4;
			end if;
		
		when S5 =>
			selector <= '0';
			En0 <= '1';
			En1 <= '1';
			dir0 <= '0';
			dir1 <= '1';
			if cont = 133 then --Contamos hasta 15
				esiguiente<=S6;
			else
				esiguiente<=S5;
			end if;
	
		when S6 =>
			selector <= '0';
			En0 <= '1';
			En1 <= '0';
			dir0 <= '0';
			dir1 <= '1';
			if cont = 250 then --Contamos hasta 15
				esiguiente<=S7;
			else
				esiguiente<=S6;
			end if;

		when S7 =>
			selector <= '0';
			En0 <= '1';
			En1 <= '1';
			dir0 <= '0';
			dir1 <= '0';
			if cont = 133 then --Contamos hasta 15
				esiguiente<=S8;
			else
				esiguiente<=S7;
			end if;

		when S8 =>
			selector <= '0';
			En0 <= '0';
			En1 <= '1';
			dir0 <= '0';
			dir1 <= '0';
			if cont = 250 then --Contamos hasta 15
				esiguiente<=S9;
			else
				esiguiente<=S8;
			end if;	

		when S9 =>
			selector <= '0';
			En0 <= '1';
			En1 <= '1';
			dir0 <= '1';
			dir1 <= '0';
			if cont = 133 then --Contamos hasta 15
				esiguiente<=S0;
			else
				esiguiente<=S9;
			end if;	
	
	end case;
end process;
	
end Behavioral;